module main

import repl

fn main() {
	println('vmonkey REPL')

	repl.start()
}
