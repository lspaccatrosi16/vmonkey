module parser

fn test_parser() {}
